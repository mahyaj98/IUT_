** Profile: "SCHEMATIC1-THIS"  [ d:\dc_rl-schematic1-this.sim ] 

** Creating circuit file "dc_rl-schematic1-this.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\dc_rl-SCHEMATIC1.net" 


.END
