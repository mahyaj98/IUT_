** Profile: "SCHEMATIC1-new"  [ D:\DC_RESISTOR\new-SCHEMATIC1-new.sim ] 

** Creating circuit file "new-SCHEMATIC1-new.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\new-SCHEMATIC1.net" 


.END
