** Profile: "SCHEMATIC1-RC"  [ D:\rc-SCHEMATIC1-RC.sim ] 

** Creating circuit file "rc-SCHEMATIC1-RC.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 2 0 1
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\rc-SCHEMATIC1.net" 


.END
